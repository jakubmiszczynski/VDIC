/*
 Copyright 2013 Ray Salemi

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at

 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 
 Last modification: 2024-10-22 AGH RSz
 */
module tpgen(fifomult_bfm bfm);
    
import fifomult_tb_pkg::*;




initial begin : tpgen
	parameter A = 100;
	parameter fifo_break = 100;
	parameter M = 100;
	bfm.reset_fifomult();

	// Corners test, parity test
	repeat (A) begin
	    begin
		    bfm.send_data();
	    end
	end
	
	repeat (fifo_break) begin
	    begin
		    bfm.send_nothing();
	    end
	end
	// Busy test
	repeat (M) begin
	    begin
		    bfm.send_data_busy_test();  
	    end
	end
	repeat (fifo_break) begin
	    begin
		    bfm.send_nothing();
	    end
	end
    $finish;
end : tpgen

endmodule : tpgen
